/*************************************************************************
 > Copyright (C) 2021 Sangfor Ltd. All rights reserved.
 > File Name   : router_defines.sv
 > Author      : bhyou
 > Mail        : bhyou@foxmail.com 
 > Created Time: Mon 19 Jul 2021 02:03:57 PM CST
 ************************************************************************/
`define SOF  2'b10
`define DATA 2'b00
`define EOF  2'b01
 
`define DataPacketSize 5
//`define DataPacketSize 35